library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use std.env.finish;

library osvvm;
use osvvm.RandomPkg.all;
use osvvm.CoveragePkg.all;

use work.DataStructures.all;

-- enter your code below
entity alu_tb is 

end alu_tb;

architecture tb of alu_tb is 
begin 

end tb;